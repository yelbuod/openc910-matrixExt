module ct_mat_idu_top (
    input         id_inst0_m_inst_vld,
    input         id_inst1_m_inst_vld,
    input         id_inst2_m_inst_vld,
    input  [22:0] id_inst0_m_data    ,
    input  [22:0] id_inst1_m_data    ,
    input  [22:0] id_inst2_m_data    ,
    output        mat_idu_stall
);



endmodule : ct_mat_idu_top